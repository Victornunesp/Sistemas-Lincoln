entity CLA_4b is
	port();
end CLA_4b;

architecture mega_soma of CLA_4b is
begin

end mega_soma;